** sch_path: /home/nwells/xschem/6_bit_flash/schematics/decoder_top.sch
**.subckt decoder_top VDD OUT5,OUT4,OUT3,OUT2,OUT1,OUT0 VSS
*+ decode_in62,decode_in61,decode_in60,decode_in59,decode_in58,decode_in57,decode_in56,decode_in55,decode_in54,decode_in53,decode_in52,decode_in51,decode_in50,decode_in49,decode_in48,decode_in47,decode_in46,decode_in45,decode_in44,decode_in43,decode_in42,decode_in41,decode_in40,decode_in39,decode_in38,decode_in37,decode_in36,decode_in35,decode_in34,decode_in33,decode_in32,decode_in31,decode_in30,decode_in29,decode_in28,decode_in27,decode_in26,decode_in25,decode_in24,decode_in23,decode_in22,decode_in21,decode_in20,decode_in19,decode_in18,decode_in17,decode_in16,decode_in15,decode_in14,decode_in13,decode_in12,decode_in11,decode_in10,decode_in9,decode_in8,decode_in7,decode_in6,decode_in5,decode_in4,decode_in3,decode_in2,decode_in1,decode_in0
*.ipin
*+ decode_in62,decode_in61,decode_in60,decode_in59,decode_in58,decode_in57,decode_in56,decode_in55,decode_in54,decode_in53,decode_in52,decode_in51,decode_in50,decode_in49,decode_in48,decode_in47,decode_in46,decode_in45,decode_in44,decode_in43,decode_in42,decode_in41,decode_in40,decode_in39,decode_in38,decode_in37,decode_in36,decode_in35,decode_in34,decode_in33,decode_in32,decode_in31,decode_in30,decode_in29,decode_in28,decode_in27,decode_in26,decode_in25,decode_in24,decode_in23,decode_in22,decode_in21,decode_in20,decode_in19,decode_in18,decode_in17,decode_in16,decode_in15,decode_in14,decode_in13,decode_in12,decode_in11,decode_in10,decode_in9,decode_in8,decode_in7,decode_in6,decode_in5,decode_in4,decode_in3,decode_in2,decode_in1,decode_in0
*.ipin VDD
*.ipin VSS
*.opin OUT5,OUT4,OUT3,OUT2,OUT1,OUT0
XR1[63] net1[63] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[62] net1[62] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[61] net1[61] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[60] net1[60] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[59] net1[59] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[58] net1[58] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[57] net1[57] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[56] net1[56] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[55] net1[55] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[54] net1[54] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[53] net1[53] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[52] net1[52] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[51] net1[51] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[50] net1[50] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[49] net1[49] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[48] net1[48] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[47] net1[47] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[46] net1[46] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[45] net1[45] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[44] net1[44] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[43] net1[43] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[42] net1[42] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[41] net1[41] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[40] net1[40] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[39] net1[39] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[38] net1[38] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[37] net1[37] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[36] net1[36] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[35] net1[35] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[34] net1[34] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[33] net1[33] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[32] net1[32] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[31] net1[31] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[30] net1[30] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[29] net1[29] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[28] net1[28] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[27] net1[27] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[26] net1[26] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[25] net1[25] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[24] net1[24] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[23] net1[23] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[22] net1[22] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[21] net1[21] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[20] net1[20] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[19] net1[19] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[18] net1[18] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[17] net1[17] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[16] net1[16] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[15] net1[15] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[14] net1[14] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[13] net1[13] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[12] net1[12] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[11] net1[11] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[10] net1[10] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[9] net1[9] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[8] net1[8] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[7] net1[7] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[6] net1[6] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[5] net1[5] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[4] net1[4] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[3] net1[3] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[2] net1[2] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[1] net1[1] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1[0] net1[0] OUT5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[63] net1[63] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[62] net1[62] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[61] net1[61] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[60] net1[60] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[59] net1[59] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[58] net1[58] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[57] net1[57] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[56] net1[56] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[55] net1[55] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[54] net1[54] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[53] net1[53] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[52] net1[52] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[51] net1[51] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[50] net1[50] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[49] net1[49] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[48] net1[48] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[47] net1[47] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[46] net1[46] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[45] net1[45] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[44] net1[44] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[43] net1[43] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[42] net1[42] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[41] net1[41] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[40] net1[40] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[39] net1[39] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[38] net1[38] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[37] net1[37] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[36] net1[36] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[35] net1[35] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[34] net1[34] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[33] net1[33] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[32] net1[32] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[31] net1[31] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[30] net1[30] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[29] net1[29] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[28] net1[28] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[27] net1[27] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[26] net1[26] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[25] net1[25] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[24] net1[24] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[23] net1[23] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[22] net1[22] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[21] net1[21] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[20] net1[20] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[19] net1[19] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[18] net1[18] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[17] net1[17] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[16] net1[16] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[15] net1[15] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[14] net1[14] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[13] net1[13] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[12] net1[12] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[11] net1[11] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[10] net1[10] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[9] net1[9] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[8] net1[8] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[7] net1[7] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[6] net1[6] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[5] net1[5] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[4] net1[4] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[3] net1[3] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[2] net1[2] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[1] net1[1] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2[0] net1[0] OUT4 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[63] net1[63] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[62] net1[62] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[61] net1[61] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[60] net1[60] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[59] net1[59] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[58] net1[58] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[57] net1[57] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[56] net1[56] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[55] net1[55] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[54] net1[54] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[53] net1[53] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[52] net1[52] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[51] net1[51] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[50] net1[50] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[49] net1[49] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[48] net1[48] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[47] net1[47] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[46] net1[46] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[45] net1[45] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[44] net1[44] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[43] net1[43] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[42] net1[42] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[41] net1[41] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[40] net1[40] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[39] net1[39] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[38] net1[38] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[37] net1[37] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[36] net1[36] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[35] net1[35] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[34] net1[34] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[33] net1[33] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[32] net1[32] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[31] net1[31] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[30] net1[30] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[29] net1[29] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[28] net1[28] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[27] net1[27] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[26] net1[26] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[25] net1[25] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[24] net1[24] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[23] net1[23] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[22] net1[22] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[21] net1[21] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[20] net1[20] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[19] net1[19] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[18] net1[18] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[17] net1[17] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[16] net1[16] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[15] net1[15] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[14] net1[14] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[13] net1[13] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[12] net1[12] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[11] net1[11] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[10] net1[10] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[9] net1[9] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[8] net1[8] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[7] net1[7] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[6] net1[6] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[5] net1[5] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[4] net1[4] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[3] net1[3] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[2] net1[2] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[1] net1[1] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3[0] net1[0] OUT3 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[63] net2[63] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[62] net2[62] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[61] net2[61] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[60] net2[60] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[59] net2[59] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[58] net2[58] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[57] net2[57] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[56] net2[56] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[55] net2[55] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[54] net2[54] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[53] net2[53] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[52] net2[52] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[51] net2[51] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[50] net2[50] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[49] net2[49] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[48] net2[48] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[47] net2[47] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[46] net2[46] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[45] net2[45] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[44] net2[44] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[43] net2[43] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[42] net2[42] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[41] net2[41] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[40] net2[40] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[39] net2[39] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[38] net2[38] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[37] net2[37] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[36] net2[36] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[35] net2[35] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[34] net2[34] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[33] net2[33] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[32] net2[32] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[31] net2[31] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[30] net2[30] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[29] net2[29] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[28] net2[28] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[27] net2[27] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[26] net2[26] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[25] net2[25] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[24] net2[24] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[23] net2[23] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[22] net2[22] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[21] net2[21] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[20] net2[20] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[19] net2[19] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[18] net2[18] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[17] net2[17] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[16] net2[16] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[15] net2[15] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[14] net2[14] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[13] net2[13] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[12] net2[12] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[11] net2[11] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[10] net2[10] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[9] net2[9] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[8] net2[8] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[7] net2[7] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[6] net2[6] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[5] net2[5] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[4] net2[4] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[3] net2[3] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[2] net2[2] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[1] net2[1] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4[0] net2[0] OUT2 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[63] net2[63] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[62] net2[62] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[61] net2[61] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[60] net2[60] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[59] net2[59] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[58] net2[58] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[57] net2[57] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[56] net2[56] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[55] net2[55] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[54] net2[54] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[53] net2[53] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[52] net2[52] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[51] net2[51] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[50] net2[50] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[49] net2[49] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[48] net2[48] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[47] net2[47] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[46] net2[46] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[45] net2[45] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[44] net2[44] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[43] net2[43] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[42] net2[42] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[41] net2[41] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[40] net2[40] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[39] net2[39] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[38] net2[38] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[37] net2[37] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[36] net2[36] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[35] net2[35] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[34] net2[34] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[33] net2[33] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[32] net2[32] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[31] net2[31] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[30] net2[30] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[29] net2[29] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[28] net2[28] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[27] net2[27] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[26] net2[26] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[25] net2[25] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[24] net2[24] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[23] net2[23] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[22] net2[22] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[21] net2[21] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[20] net2[20] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[19] net2[19] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[18] net2[18] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[17] net2[17] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[16] net2[16] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[15] net2[15] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[14] net2[14] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[13] net2[13] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[12] net2[12] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[11] net2[11] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[10] net2[10] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[9] net2[9] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[8] net2[8] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[7] net2[7] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[6] net2[6] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[5] net2[5] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[4] net2[4] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[3] net2[3] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[2] net2[2] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[1] net2[1] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5[0] net2[0] OUT1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[63] net2[63] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[62] net2[62] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[61] net2[61] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[60] net2[60] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[59] net2[59] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[58] net2[58] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[57] net2[57] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[56] net2[56] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[55] net2[55] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[54] net2[54] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[53] net2[53] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[52] net2[52] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[51] net2[51] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[50] net2[50] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[49] net2[49] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[48] net2[48] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[47] net2[47] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[46] net2[46] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[45] net2[45] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[44] net2[44] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[43] net2[43] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[42] net2[42] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[41] net2[41] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[40] net2[40] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[39] net2[39] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[38] net2[38] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[37] net2[37] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[36] net2[36] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[35] net2[35] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[34] net2[34] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[33] net2[33] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[32] net2[32] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[31] net2[31] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[30] net2[30] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[29] net2[29] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[28] net2[28] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[27] net2[27] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[26] net2[26] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[25] net2[25] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[24] net2[24] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[23] net2[23] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[22] net2[22] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[21] net2[21] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[20] net2[20] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[19] net2[19] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[18] net2[18] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[17] net2[17] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[16] net2[16] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[15] net2[15] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[14] net2[14] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[13] net2[13] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[12] net2[12] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[11] net2[11] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[10] net2[10] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[9] net2[9] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[8] net2[8] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[7] net2[7] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[6] net2[6] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[5] net2[5] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[4] net2[4] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[3] net2[3] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[2] net2[2] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[1] net2[1] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6[0] net2[0] OUT0 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
**.ends
.end
