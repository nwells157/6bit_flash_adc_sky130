** sch_path: /home/nwells/xschem/6_bit_flash/schematics/comp_top.sch
**.subckt comp_top VDD
*+ vout62,vout61,vout60,vout59,vout58,vout57,vout56,vout55,vout54,vout53,vout52,vout51,vout50,vout49,vout48,vout47,vout46,vout45,vout44,vout43,vout42,vout41,vout40,vout39,vout38,vout37,vout36,vout35,vout34,vout33,vout32,vout31,vout30,vout29,vout28,vout27,vout26,vout25,vout24,vout23,vout22,vout21,vout20,vout19,vout18,vout17,vout16,vout15,vout14,vout13,vout12,vout11,vout10,vout9,vout8,vout7,vout6,vout5,vout4,vout3,vout2,vout1,vout0 VSS
*+ vref62,vref61,vref60,vref59,vref58,vref57,vref56,vref55,vref54,vref53,vref52,vref51,vref50,vref49,vref48,vref47,vref46,vref45,vref44,vref43,vref42,vref41,vref40,vref39,vref38,vref37,vref36,vref35,vref34,vref33,vref32,vref31,vref30,vref29,vref28,vref27,vref26,vref25,vref24,vref23,vref22,vref21,vref20,vref19,vref18,vref17,vref16,vref15,vref14,vref13,vref12,vref11,vref10,vref9,vref8,vref7,vref6,vref5,vref4,vref3,vref2,vref1,vref0 VIN clk
*.opin
*+ vout62,vout61,vout60,vout59,vout58,vout57,vout56,vout55,vout54,vout53,vout52,vout51,vout50,vout49,vout48,vout47,vout46,vout45,vout44,vout43,vout42,vout41,vout40,vout39,vout38,vout37,vout36,vout35,vout34,vout33,vout32,vout31,vout30,vout29,vout28,vout27,vout26,vout25,vout24,vout23,vout22,vout21,vout20,vout19,vout18,vout17,vout16,vout15,vout14,vout13,vout12,vout11,vout10,vout9,vout8,vout7,vout6,vout5,vout4,vout3,vout2,vout1,vout0
*.ipin VDD
*.ipin VSS
*.ipin
*+ vref62,vref61,vref60,vref59,vref58,vref57,vref56,vref55,vref54,vref53,vref52,vref51,vref50,vref49,vref48,vref47,vref46,vref45,vref44,vref43,vref42,vref41,vref40,vref39,vref38,vref37,vref36,vref35,vref34,vref33,vref32,vref31,vref30,vref29,vref28,vref27,vref26,vref25,vref24,vref23,vref22,vref21,vref20,vref19,vref18,vref17,vref16,vref15,vref14,vref13,vref12,vref11,vref10,vref9,vref8,vref7,vref6,vref5,vref4,vref3,vref2,vref1,vref0
*.ipin VIN
*.ipin clk
xCOMP62 vout62 VDD VSS VIN vref62 clk comp
xCOMP61 vout61 VDD VSS VIN vref61 clk comp
xCOMP60 vout60 VDD VSS VIN vref60 clk comp
xCOMP59 vout59 VDD VSS VIN vref59 clk comp
xCOMP58 vout58 VDD VSS VIN vref58 clk comp
xCOMP57 vout57 VDD VSS VIN vref57 clk comp
xCOMP56 vout56 VDD VSS VIN vref56 clk comp
xCOMP55 vout55 VDD VSS VIN vref55 clk comp
xCOMP54 vout54 VDD VSS VIN vref54 clk comp
xCOMP53 vout53 VDD VSS VIN vref53 clk comp
xCOMP52 vout52 VDD VSS VIN vref52 clk comp
xCOMP51 vout51 VDD VSS VIN vref51 clk comp
xCOMP50 vout50 VDD VSS VIN vref50 clk comp
xCOMP49 vout49 VDD VSS VIN vref49 clk comp
xCOMP48 vout48 VDD VSS VIN vref48 clk comp
xCOMP47 vout47 VDD VSS VIN vref47 clk comp
xCOMP46 vout46 VDD VSS VIN vref46 clk comp
xCOMP45 vout45 VDD VSS VIN vref45 clk comp
xCOMP44 vout44 VDD VSS VIN vref44 clk comp
xCOMP43 vout43 VDD VSS VIN vref43 clk comp
xCOMP42 vout42 VDD VSS VIN vref42 clk comp
xCOMP41 vout41 VDD VSS VIN vref41 clk comp
xCOMP40 vout40 VDD VSS VIN vref40 clk comp
xCOMP39 vout39 VDD VSS VIN vref39 clk comp
xCOMP38 vout38 VDD VSS VIN vref38 clk comp
xCOMP37 vout37 VDD VSS VIN vref37 clk comp
xCOMP36 vout36 VDD VSS VIN vref36 clk comp
xCOMP35 vout35 VDD VSS VIN vref35 clk comp
xCOMP34 vout34 VDD VSS VIN vref34 clk comp
xCOMP33 vout33 VDD VSS VIN vref33 clk comp
xCOMP32 vout32 VDD VSS VIN vref32 clk comp
xCOMP31 vout31 VDD VSS VIN vref31 clk comp
xCOMP30 vout30 VDD VSS VIN vref30 clk comp
xCOMP29 vout29 VDD VSS VIN vref29 clk comp
xCOMP28 vout28 VDD VSS VIN vref28 clk comp
xCOMP27 vout27 VDD VSS VIN vref27 clk comp
xCOMP26 vout26 VDD VSS VIN vref26 clk comp
xCOMP25 vout25 VDD VSS VIN vref25 clk comp
xCOMP24 vout24 VDD VSS VIN vref24 clk comp
xCOMP23 vout23 VDD VSS VIN vref23 clk comp
xCOMP22 vout22 VDD VSS VIN vref22 clk comp
xCOMP21 vout21 VDD VSS VIN vref21 clk comp
xCOMP20 vout20 VDD VSS VIN vref20 clk comp
xCOMP19 vout19 VDD VSS VIN vref19 clk comp
xCOMP18 vout18 VDD VSS VIN vref18 clk comp
xCOMP17 vout17 VDD VSS VIN vref17 clk comp
xCOMP16 vout16 VDD VSS VIN vref16 clk comp
xCOMP15 vout15 VDD VSS VIN vref15 clk comp
xCOMP14 vout14 VDD VSS VIN vref14 clk comp
xCOMP13 vout13 VDD VSS VIN vref13 clk comp
xCOMP12 vout12 VDD VSS VIN vref12 clk comp
xCOMP11 vout11 VDD VSS VIN vref11 clk comp
xCOMP10 vout10 VDD VSS VIN vref10 clk comp
xCOMP9 vout9 VDD VSS VIN vref9 clk comp
xCOMP8 vout8 VDD VSS VIN vref8 clk comp
xCOMP7 vout7 VDD VSS VIN vref7 clk comp
xCOMP6 vout6 VDD VSS VIN vref6 clk comp
xCOMP5 vout5 VDD VSS VIN vref5 clk comp
xCOMP4 vout4 VDD VSS VIN vref4 clk comp
xCOMP3 vout3 VDD VSS VIN vref3 clk comp
xCOMP2 vout2 VDD VSS VIN vref2 clk comp
xCOMP1 vout1 VDD VSS VIN vref1 clk comp
xCOMP0 vout0 VDD VSS VIN vref0 clk comp
**.ends

* expanding   symbol:  schematics/comp.sym # of pins=6
** sym_path: /home/nwells/xschem/6_bit_flash/schematics/comp.sym
** sch_path: /home/nwells/xschem/6_bit_flash/schematics/comp.sch
.subckt comp vout vdd vss vinp vinn clk
*.ipin vdd
*.opin vout
*.ipin vss
*.ipin vinp
*.ipin vinn
*.ipin clk
XM1 vinp_d vinp vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM2 vinn_d vinn vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM3 voutn voutp vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=7.5 nf=1 ad=2.175 as=2.175 pd=15.58 ps=15.58 nrd=0.0386666666666667
+ nrs=0.0386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM4 voutp voutn vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=7.5 nf=1 ad=2.175 as=2.175 pd=15.58 ps=15.58 nrd=0.0386666666666667
+ nrs=0.0386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM5 vinp_d vinn_d vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=7.5 nf=1 ad=2.175 as=2.175 pd=15.58 ps=15.58 nrd=0.0386666666666667
+ nrs=0.0386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM6 vinn_d vinp_d vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=7.5 nf=1 ad=2.175 as=2.175 pd=15.58 ps=15.58 nrd=0.0386666666666667
+ nrs=0.0386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM7 voutn clk vinp_d vss sky130_fd_pr__nfet_01v8 L=0.18 W=1.5 nf=1 ad=0.435 as=0.435 pd=3.58 ps=3.58 nrd=0.193333333333333
+ nrs=0.193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM8 voutp clk vinn_d vss sky130_fd_pr__nfet_01v8 L=0.18 W=1.5 nf=1 ad=0.435 as=0.435 pd=3.58 ps=3.58 nrd=0.193333333333333
+ nrs=0.193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM9 voutn clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=4 nf=1 ad=1.16 as=1.16 pd=8.58 ps=8.58 nrd=0.0725 nrs=0.0725 sa=0 sb=0 sd=0
+ mult=1 m=1
XM10 voutp clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=4 nf=1 ad=1.16 as=1.16 pd=8.58 ps=8.58 nrd=0.0725 nrs=0.0725 sa=0 sb=0
+ sd=0 mult=1 m=1
xBUFF voutp vss vss vdd vdd voutp_buff sky130_fd_sc_hd__buf_6
xBUFF1 voutn vss vss vdd vdd voutn_buff sky130_fd_sc_hd__buf_6
I0 pa_m1_s vss 10u
XM11 v_m1_d voutp_buff pa_m1_s vss sky130_fd_pr__nfet_01v8 L=0.15 W=50 nf=1 ad=14.5 as=14.5 pd=100.58 ps=100.58 nrd=0.0058
+ nrs=0.0058 sa=0 sb=0 sd=0 mult=1 m=1
XM12 vout voutn_buff pa_m1_s vss sky130_fd_pr__nfet_01v8 L=0.15 W=50 nf=1 ad=14.5 as=14.5 pd=100.58 ps=100.58 nrd=0.0058
+ nrs=0.0058 sa=0 sb=0 sd=0 mult=1 m=1
XM13 v_m1_d v_m1_d vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0
+ sd=0 mult=1 m=1
XM14 vout v_m1_d vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
.ends

.end
