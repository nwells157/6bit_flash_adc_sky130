** sch_path: /home/nwells/xschem/6_bit_flash/schematics/ideal_decoder_2bit.sch
**.subckt ideal_decoder_2bit out1,out0 vdd vss vref in3,in2,in1,in0
*.ipin vdd
*.ipin vss
*.ipin vref
*.ipin in3,in2,in1,in0
*.opin out1,out0
**.ends
.end
