** sch_path: /home/nwells/xschem/6_bit_flash/schematics/adc_top.sch
**.subckt adc_top OUT5,OUT4,OUT3,OUT2,OUT1,OUT0 VDD
*+ vref62,vref61,vref60,vref59,vref58,vref57,vref56,vref55,vref54,vref53,vref52,vref51,vref50,vref49,vref48,vref47,vref46,vref45,vref44,vref43,vref42,vref41,vref40,vref39,vref38,vref37,vref36,vref35,vref34,vref33,vref32,vref31,vref30,vref29,vref28,vref27,vref26,vref25,vref24,vref23,vref22,vref21,vref20,vref19,vref18,vref17,vref16,vref15,vref14,vref13,vref12,vref11,vref10,vref9,vref8,vref7,vref6,vref5,vref4,vref3,vref2,vref1,vref0 VSS
*+ comp_out62,comp_out61,comp_out60,comp_out59,comp_out58,comp_out57,comp_out56,comp_out55,comp_out54,comp_out53,comp_out52,comp_out51,comp_out50,comp_out49,comp_out48,comp_out47,comp_out46,comp_out45,comp_out44,comp_out43,comp_out42,comp_out41,comp_out40,comp_out39,comp_out38,comp_out37,comp_out36,comp_out35,comp_out34,comp_out33,comp_out32,comp_out31,comp_out30,comp_out29,comp_out28,comp_out27,comp_out26,comp_out25,comp_out24,comp_out23,comp_out22,comp_out21,comp_out20,comp_out19,comp_out18,comp_out17,comp_out16,comp_out15,comp_out14,comp_out13,comp_out12,comp_out11,comp_out10,comp_out9,comp_out8,comp_out7,comp_out6,comp_out5,comp_out4,comp_out3,comp_out2,comp_out1,comp_out0 VIN VREF clk
*.ipin VDD
*.ipin VSS
*.ipin VIN
*.ipin VREF
*.opin OUT5,OUT4,OUT3,OUT2,OUT1,OUT0
*.iopin
*+ vref62,vref61,vref60,vref59,vref58,vref57,vref56,vref55,vref54,vref53,vref52,vref51,vref50,vref49,vref48,vref47,vref46,vref45,vref44,vref43,vref42,vref41,vref40,vref39,vref38,vref37,vref36,vref35,vref34,vref33,vref32,vref31,vref30,vref29,vref28,vref27,vref26,vref25,vref24,vref23,vref22,vref21,vref20,vref19,vref18,vref17,vref16,vref15,vref14,vref13,vref12,vref11,vref10,vref9,vref8,vref7,vref6,vref5,vref4,vref3,vref2,vref1,vref0
*.iopin
*+ comp_out62,comp_out61,comp_out60,comp_out59,comp_out58,comp_out57,comp_out56,comp_out55,comp_out54,comp_out53,comp_out52,comp_out51,comp_out50,comp_out49,comp_out48,comp_out47,comp_out46,comp_out45,comp_out44,comp_out43,comp_out42,comp_out41,comp_out40,comp_out39,comp_out38,comp_out37,comp_out36,comp_out35,comp_out34,comp_out33,comp_out32,comp_out31,comp_out30,comp_out29,comp_out28,comp_out27,comp_out26,comp_out25,comp_out24,comp_out23,comp_out22,comp_out21,comp_out20,comp_out19,comp_out18,comp_out17,comp_out16,comp_out15,comp_out14,comp_out13,comp_out12,comp_out11,comp_out10,comp_out9,comp_out8,comp_out7,comp_out6,comp_out5,comp_out4,comp_out3,comp_out2,comp_out1,comp_out0
*.ipin clk
xREF_LADDER VDD vref62 vref61 vref60 vref59 vref58 vref57 vref56 vref55 vref54 vref53 vref52 vref51 vref50 vref49 vref48 vref47
+ vref46 vref45 vref44 vref43 vref42 vref41 vref40 vref39 vref38 vref37 vref36 vref35 vref34 vref33 vref32 vref31 vref30 vref29 vref28
+ vref27 vref26 vref25 vref24 vref23 vref22 vref21 vref20 vref19 vref18 vref17 vref16 vref15 vref14 vref13 vref12 vref11 vref10 vref9
+ vref8 vref7 vref6 vref5 vref4 vref3 vref2 vref1 vref0 VSS ref_ladder_top
xDECODER_6BIT_VERILOGA VDD OUT5 OUT4 OUT3 OUT2 OUT1 OUT0 comp_out62 comp_out61 comp_out60 comp_out59 comp_out58 comp_out57
+ comp_out56 comp_out55 comp_out54 comp_out53 comp_out52 comp_out51 comp_out50 comp_out49 comp_out48 comp_out47 comp_out46 comp_out45
+ comp_out44 comp_out43 comp_out42 comp_out41 comp_out40 comp_out39 comp_out38 comp_out37 comp_out36 comp_out35 comp_out34 comp_out33
+ comp_out32 comp_out31 comp_out30 comp_out29 comp_out28 comp_out27 comp_out26 comp_out25 comp_out24 comp_out23 comp_out22 comp_out21
+ comp_out20 comp_out19 comp_out18 comp_out17 comp_out16 comp_out15 comp_out14 comp_out13 comp_out12 comp_out11 comp_out10 comp_out9 comp_out8
+ comp_out7 comp_out6 comp_out5 comp_out4 comp_out3 comp_out2 comp_out1 comp_out0 VSS VREF decoder_6bit_cell
xCOMP_TOP VDD comp_out62 comp_out61 comp_out60 comp_out59 comp_out58 comp_out57 comp_out56 comp_out55 comp_out54 comp_out53
+ comp_out52 comp_out51 comp_out50 comp_out49 comp_out48 comp_out47 comp_out46 comp_out45 comp_out44 comp_out43 comp_out42 comp_out41
+ comp_out40 comp_out39 comp_out38 comp_out37 comp_out36 comp_out35 comp_out34 comp_out33 comp_out32 comp_out31 comp_out30 comp_out29
+ comp_out28 comp_out27 comp_out26 comp_out25 comp_out24 comp_out23 comp_out22 comp_out21 comp_out20 comp_out19 comp_out18 comp_out17
+ comp_out16 comp_out15 comp_out14 comp_out13 comp_out12 comp_out11 comp_out10 comp_out9 comp_out8 comp_out7 comp_out6 comp_out5 comp_out4
+ comp_out3 comp_out2 comp_out1 comp_out0 VSS vref62 vref61 vref60 vref59 vref58 vref57 vref56 vref55 vref54 vref53 vref52 vref51 vref50
+ vref49 vref48 vref47 vref46 vref45 vref44 vref43 vref42 vref41 vref40 vref39 vref38 vref37 vref36 vref35 vref34 vref33 vref32 vref31
+ vref30 vref29 vref28 vref27 vref26 vref25 vref24 vref23 vref22 vref21 vref20 vref19 vref18 vref17 vref16 vref15 vref14 vref13 vref12
+ vref11 vref10 vref9 vref8 vref7 vref6 vref5 vref4 vref3 vref2 vref1 vref0 VIN clk comp_top
**.ends

* expanding   symbol:  schematics/ref_ladder_top.sym # of pins=3
** sym_path: /home/nwells/xschem/6_bit_flash/schematics/ref_ladder_top.sym
** sch_path: /home/nwells/xschem/6_bit_flash/schematics/ref_ladder_top.sch
.subckt ref_ladder_top VDD vref62 vref61 vref60 vref59 vref58 vref57 vref56 vref55 vref54 vref53 vref52 vref51 vref50 vref49
+ vref48 vref47 vref46 vref45 vref44 vref43 vref42 vref41 vref40 vref39 vref38 vref37 vref36 vref35 vref34 vref33 vref32 vref31 vref30
+ vref29 vref28 vref27 vref26 vref25 vref24 vref23 vref22 vref21 vref20 vref19 vref18 vref17 vref16 vref15 vref14 vref13 vref12 vref11
+ vref10 vref9 vref8 vref7 vref6 vref5 vref4 vref3 vref2 vref1 vref0 VSS
*.ipin VDD
*.opin
*+ vref62,vref61,vref60,vref59,vref58,vref57,vref56,vref55,vref54,vref53,vref52,vref51,vref50,vref49,vref48,vref47,vref46,vref45,vref44,vref43,vref42,vref41,vref40,vref39,vref38,vref37,vref36,vref35,vref34,vref33,vref32,vref31,vref30,vref29,vref28,vref27,vref26,vref25,vref24,vref23,vref22,vref21,vref20,vref19,vref18,vref17,vref16,vref15,vref14,vref13,vref12,vref11,vref10,vref9,vref8,vref7,vref6,vref5,vref4,vref3,vref2,vref1,vref0
*.ipin VSS
XR1[63] vref62 VDD VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[62] vref61 vref62 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[61] vref60 vref61 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[60] vref59 vref60 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[59] vref58 vref59 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[58] vref57 vref58 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[57] vref56 vref57 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[56] vref55 vref56 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[55] vref54 vref55 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[54] vref53 vref54 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[53] vref52 vref53 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[52] vref51 vref52 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[51] vref50 vref51 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[50] vref49 vref50 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[49] vref48 vref49 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[48] vref47 vref48 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[47] vref46 vref47 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[46] vref45 vref46 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[45] vref44 vref45 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[44] vref43 vref44 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[43] vref42 vref43 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[42] vref41 vref42 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[41] vref40 vref41 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[40] vref39 vref40 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[39] vref38 vref39 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[38] vref37 vref38 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[37] vref36 vref37 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[36] vref35 vref36 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[35] vref34 vref35 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[34] vref33 vref34 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[33] vref32 vref33 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[32] vref31 vref32 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[31] vref30 vref31 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[30] vref29 vref30 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[29] vref28 vref29 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[28] vref27 vref28 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[27] vref26 vref27 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[26] vref25 vref26 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[25] vref24 vref25 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[24] vref23 vref24 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[23] vref22 vref23 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[22] vref21 vref22 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[21] vref20 vref21 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[20] vref19 vref20 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[19] vref18 vref19 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[18] vref17 vref18 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[17] vref16 vref17 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[16] vref15 vref16 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[15] vref14 vref15 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[14] vref13 vref14 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[13] vref12 vref13 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[12] vref11 vref12 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[11] vref10 vref11 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[10] vref9 vref10 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[9] vref8 vref9 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[8] vref7 vref8 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[7] vref6 vref7 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[6] vref5 vref6 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[5] vref4 vref5 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[4] vref3 vref4 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[3] vref2 vref3 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[2] vref1 vref2 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[1] vref0 vref1 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
XR1[0] VSS vref0 VSS sky130_fd_pr__res_high_po W=7 L=1 mult=1 m=1
.ends


* expanding   symbol:  schematics/comp_top_ideal.sym # of pins=5
** sym_path: /home/nwells/xschem/6_bit_flash/schematics/comp_top_ideal.sym
** sch_path: /home/nwells/xschem/6_bit_flash/schematics/comp_top_ideal.sch
.subckt comp_top_ideal vout62 vout61 vout60 vout59 vout58 vout57 vout56 vout55 vout54 vout53 vout52 vout51 vout50 vout49 vout48
+ vout47 vout46 vout45 vout44 vout43 vout42 vout41 vout40 vout39 vout38 vout37 vout36 vout35 vout34 vout33 vout32 vout31 vout30 vout29
+ vout28 vout27 vout26 vout25 vout24 vout23 vout22 vout21 vout20 vout19 vout18 vout17 vout16 vout15 vout14 vout13 vout12 vout11 vout10
+ vout9 vout8 vout7 vout6 vout5 vout4 vout3 vout2 vout1 vout0 VDD VSS vref62 vref61 vref60 vref59 vref58 vref57 vref56 vref55 vref54
+ vref53 vref52 vref51 vref50 vref49 vref48 vref47 vref46 vref45 vref44 vref43 vref42 vref41 vref40 vref39 vref38 vref37 vref36 vref35
+ vref34 vref33 vref32 vref31 vref30 vref29 vref28 vref27 vref26 vref25 vref24 vref23 vref22 vref21 vref20 vref19 vref18 vref17 vref16
+ vref15 vref14 vref13 vref12 vref11 vref10 vref9 vref8 vref7 vref6 vref5 vref4 vref3 vref2 vref1 vref0 VIN
*.opin
*+ vout62,vout61,vout60,vout59,vout58,vout57,vout56,vout55,vout54,vout53,vout52,vout51,vout50,vout49,vout48,vout47,vout46,vout45,vout44,vout43,vout42,vout41,vout40,vout39,vout38,vout37,vout36,vout35,vout34,vout33,vout32,vout31,vout30,vout29,vout28,vout27,vout26,vout25,vout24,vout23,vout22,vout21,vout20,vout19,vout18,vout17,vout16,vout15,vout14,vout13,vout12,vout11,vout10,vout9,vout8,vout7,vout6,vout5,vout4,vout3,vout2,vout1,vout0
*.ipin VDD
*.ipin VSS
*.ipin
*+ vref62,vref61,vref60,vref59,vref58,vref57,vref56,vref55,vref54,vref53,vref52,vref51,vref50,vref49,vref48,vref47,vref46,vref45,vref44,vref43,vref42,vref41,vref40,vref39,vref38,vref37,vref36,vref35,vref34,vref33,vref32,vref31,vref30,vref29,vref28,vref27,vref26,vref25,vref24,vref23,vref22,vref21,vref20,vref19,vref18,vref17,vref16,vref15,vref14,vref13,vref12,vref11,vref10,vref9,vref8,vref7,vref6,vref5,vref4,vref3,vref2,vref1,vref0
*.ipin VIN
xVERILOG_A_COMP62 VDD VSS VIN vref62 vout62 ideal_comp_cell
xVERILOG_A_COMP61 VDD VSS VIN vref61 vout61 ideal_comp_cell
xVERILOG_A_COMP60 VDD VSS VIN vref60 vout60 ideal_comp_cell
xVERILOG_A_COMP59 VDD VSS VIN vref59 vout59 ideal_comp_cell
xVERILOG_A_COMP58 VDD VSS VIN vref58 vout58 ideal_comp_cell
xVERILOG_A_COMP57 VDD VSS VIN vref57 vout57 ideal_comp_cell
xVERILOG_A_COMP56 VDD VSS VIN vref56 vout56 ideal_comp_cell
xVERILOG_A_COMP55 VDD VSS VIN vref55 vout55 ideal_comp_cell
xVERILOG_A_COMP54 VDD VSS VIN vref54 vout54 ideal_comp_cell
xVERILOG_A_COMP53 VDD VSS VIN vref53 vout53 ideal_comp_cell
xVERILOG_A_COMP52 VDD VSS VIN vref52 vout52 ideal_comp_cell
xVERILOG_A_COMP51 VDD VSS VIN vref51 vout51 ideal_comp_cell
xVERILOG_A_COMP50 VDD VSS VIN vref50 vout50 ideal_comp_cell
xVERILOG_A_COMP49 VDD VSS VIN vref49 vout49 ideal_comp_cell
xVERILOG_A_COMP48 VDD VSS VIN vref48 vout48 ideal_comp_cell
xVERILOG_A_COMP47 VDD VSS VIN vref47 vout47 ideal_comp_cell
xVERILOG_A_COMP46 VDD VSS VIN vref46 vout46 ideal_comp_cell
xVERILOG_A_COMP45 VDD VSS VIN vref45 vout45 ideal_comp_cell
xVERILOG_A_COMP44 VDD VSS VIN vref44 vout44 ideal_comp_cell
xVERILOG_A_COMP43 VDD VSS VIN vref43 vout43 ideal_comp_cell
xVERILOG_A_COMP42 VDD VSS VIN vref42 vout42 ideal_comp_cell
xVERILOG_A_COMP41 VDD VSS VIN vref41 vout41 ideal_comp_cell
xVERILOG_A_COMP40 VDD VSS VIN vref40 vout40 ideal_comp_cell
xVERILOG_A_COMP39 VDD VSS VIN vref39 vout39 ideal_comp_cell
xVERILOG_A_COMP38 VDD VSS VIN vref38 vout38 ideal_comp_cell
xVERILOG_A_COMP37 VDD VSS VIN vref37 vout37 ideal_comp_cell
xVERILOG_A_COMP36 VDD VSS VIN vref36 vout36 ideal_comp_cell
xVERILOG_A_COMP35 VDD VSS VIN vref35 vout35 ideal_comp_cell
xVERILOG_A_COMP34 VDD VSS VIN vref34 vout34 ideal_comp_cell
xVERILOG_A_COMP33 VDD VSS VIN vref33 vout33 ideal_comp_cell
xVERILOG_A_COMP32 VDD VSS VIN vref32 vout32 ideal_comp_cell
xVERILOG_A_COMP31 VDD VSS VIN vref31 vout31 ideal_comp_cell
xVERILOG_A_COMP30 VDD VSS VIN vref30 vout30 ideal_comp_cell
xVERILOG_A_COMP29 VDD VSS VIN vref29 vout29 ideal_comp_cell
xVERILOG_A_COMP28 VDD VSS VIN vref28 vout28 ideal_comp_cell
xVERILOG_A_COMP27 VDD VSS VIN vref27 vout27 ideal_comp_cell
xVERILOG_A_COMP26 VDD VSS VIN vref26 vout26 ideal_comp_cell
xVERILOG_A_COMP25 VDD VSS VIN vref25 vout25 ideal_comp_cell
xVERILOG_A_COMP24 VDD VSS VIN vref24 vout24 ideal_comp_cell
xVERILOG_A_COMP23 VDD VSS VIN vref23 vout23 ideal_comp_cell
xVERILOG_A_COMP22 VDD VSS VIN vref22 vout22 ideal_comp_cell
xVERILOG_A_COMP21 VDD VSS VIN vref21 vout21 ideal_comp_cell
xVERILOG_A_COMP20 VDD VSS VIN vref20 vout20 ideal_comp_cell
xVERILOG_A_COMP19 VDD VSS VIN vref19 vout19 ideal_comp_cell
xVERILOG_A_COMP18 VDD VSS VIN vref18 vout18 ideal_comp_cell
xVERILOG_A_COMP17 VDD VSS VIN vref17 vout17 ideal_comp_cell
xVERILOG_A_COMP16 VDD VSS VIN vref16 vout16 ideal_comp_cell
xVERILOG_A_COMP15 VDD VSS VIN vref15 vout15 ideal_comp_cell
xVERILOG_A_COMP14 VDD VSS VIN vref14 vout14 ideal_comp_cell
xVERILOG_A_COMP13 VDD VSS VIN vref13 vout13 ideal_comp_cell
xVERILOG_A_COMP12 VDD VSS VIN vref12 vout12 ideal_comp_cell
xVERILOG_A_COMP11 VDD VSS VIN vref11 vout11 ideal_comp_cell
xVERILOG_A_COMP10 VDD VSS VIN vref10 vout10 ideal_comp_cell
xVERILOG_A_COMP9 VDD VSS VIN vref9 vout9 ideal_comp_cell
xVERILOG_A_COMP8 VDD VSS VIN vref8 vout8 ideal_comp_cell
xVERILOG_A_COMP7 VDD VSS VIN vref7 vout7 ideal_comp_cell
xVERILOG_A_COMP6 VDD VSS VIN vref6 vout6 ideal_comp_cell
xVERILOG_A_COMP5 VDD VSS VIN vref5 vout5 ideal_comp_cell
xVERILOG_A_COMP4 VDD VSS VIN vref4 vout4 ideal_comp_cell
xVERILOG_A_COMP3 VDD VSS VIN vref3 vout3 ideal_comp_cell
xVERILOG_A_COMP2 VDD VSS VIN vref2 vout2 ideal_comp_cell
xVERILOG_A_COMP1 VDD VSS VIN vref1 vout1 ideal_comp_cell
xVERILOG_A_COMP0 VDD VSS VIN vref0 vout0 ideal_comp_cell
.ends


* expanding   symbol:  schematics/decoder_top.sym # of pins=4
** sym_path: /home/nwells/xschem/6_bit_flash/schematics/decoder_top.sym
** sch_path: /home/nwells/xschem/6_bit_flash/schematics/decoder_top.sch
.subckt decoder_top VDD OUT5 OUT4 OUT3 OUT2 OUT1 OUT0 VSS decode_in62 decode_in61 decode_in60 decode_in59 decode_in58 decode_in57
+ decode_in56 decode_in55 decode_in54 decode_in53 decode_in52 decode_in51 decode_in50 decode_in49 decode_in48 decode_in47 decode_in46
+ decode_in45 decode_in44 decode_in43 decode_in42 decode_in41 decode_in40 decode_in39 decode_in38 decode_in37 decode_in36 decode_in35
+ decode_in34 decode_in33 decode_in32 decode_in31 decode_in30 decode_in29 decode_in28 decode_in27 decode_in26 decode_in25 decode_in24
+ decode_in23 decode_in22 decode_in21 decode_in20 decode_in19 decode_in18 decode_in17 decode_in16 decode_in15 decode_in14 decode_in13
+ decode_in12 decode_in11 decode_in10 decode_in9 decode_in8 decode_in7 decode_in6 decode_in5 decode_in4 decode_in3 decode_in2 decode_in1
+ decode_in0
*.ipin
*+ decode_in62,decode_in61,decode_in60,decode_in59,decode_in58,decode_in57,decode_in56,decode_in55,decode_in54,decode_in53,decode_in52,decode_in51,decode_in50,decode_in49,decode_in48,decode_in47,decode_in46,decode_in45,decode_in44,decode_in43,decode_in42,decode_in41,decode_in40,decode_in39,decode_in38,decode_in37,decode_in36,decode_in35,decode_in34,decode_in33,decode_in32,decode_in31,decode_in30,decode_in29,decode_in28,decode_in27,decode_in26,decode_in25,decode_in24,decode_in23,decode_in22,decode_in21,decode_in20,decode_in19,decode_in18,decode_in17,decode_in16,decode_in15,decode_in14,decode_in13,decode_in12,decode_in11,decode_in10,decode_in9,decode_in8,decode_in7,decode_in6,decode_in5,decode_in4,decode_in3,decode_in2,decode_in1,decode_in0
*.ipin VDD
*.ipin VSS
*.opin OUT5,OUT4,OUT3,OUT2,OUT1,OUT0
xOut0 decode_in0 decode_in2 decode_in4 decode_in6 decode_in8 decode_in10 decode_in12 decode_in14 decode_in16 decode_in18
+ decode_in20 decode_in22 decode_in24 decode_in26 decode_in28 decode_in30 decode_in32 decode_in34 decode_in36 decode_in38 decode_in40
+ decode_in42 decode_in44 decode_in46 decode_in48 decode_in50 decode_in52 decode_in54 decode_in56 decode_in58 decode_in60 decode_in62 OUT0 VDD
+ VDD VSS VSS decode_in1 decode_in3 decode_in5 decode_in7 decode_in9 decode_in11 decode_in13 decode_in15 decode_in17 decode_in19
+ decode_in21 decode_in23 decode_in25 decode_in27 decode_in29 decode_in31 decode_in33 decode_in35 decode_in37 decode_in39 decode_in41
+ decode_in43 decode_in45 decode_in47 decode_in49 decode_in51 decode_in53 decode_in55 decode_in57 decode_in59 decode_in61 or_32
xOut1 decode_in1 decode_in2 decode_in5 decode_in6 decode_in9 decode_in10 decode_in13 decode_in14 decode_in17 decode_in18
+ decode_in21 decode_in22 decode_in25 decode_in26 decode_in29 decode_in30 decode_in33 decode_in34 decode_in37 decode_in38 decode_in41
+ decode_in42 decode_in45 decode_in46 decode_in49 decode_in50 decode_in53 decode_in54 decode_in57 decode_in58 decode_in61 decode_in62 OUT1 VDD
+ VDD VSS VSS decode_in2 decode_in3 decode_in6 decode_in7 decode_in10 decode_in11 decode_in14 decode_in15 decode_in18 decode_in19
+ decode_in22 decode_in23 decode_in26 decode_in27 decode_in30 decode_in31 decode_in34 decode_in35 decode_in38 decode_in39 decode_in42
+ decode_in43 decode_in46 decode_in47 decode_in50 decode_in51 decode_in54 decode_in55 decode_in58 decode_in59 decode_in62 or_32
xOut2 decode_in3 decode_in4 decode_in5 decode_in6 decode_in11 decode_in12 decode_in13 decode_in14 decode_in19 decode_in20
+ decode_in21 decode_in22 decode_in27 decode_in28 decode_in29 decode_in30 decode_in35 decode_in36 decode_in37 decode_in38 decode_in43
+ decode_in44 decode_in45 decode_in46 decode_in51 decode_in52 decode_in53 decode_in54 decode_in59 decode_in60 decode_in61 decode_in62 OUT2 VDD
+ VDD VSS VSS decode_in4 decode_in5 decode_in6 decode_in7 decode_in12 decode_in13 decode_in14 decode_in15 decode_in20 decode_in21
+ decode_in22 decode_in23 decode_in28 decode_in29 decode_in30 decode_in31 decode_in36 decode_in37 decode_in38 decode_in39 decode_in44
+ decode_in45 decode_in46 decode_in47 decode_in52 decode_in53 decode_in54 decode_in55 decode_in60 decode_in61 decode_in62 or_32
xOut3 decode_in7 decode_in8 decode_in9 decode_in10 decode_in11 decode_in12 decode_in13 decode_in14 decode_in23 decode_in24
+ decode_in25 decode_in26 decode_in27 decode_in28 decode_in29 decode_in30 decode_in39 decode_in40 decode_in41 decode_in42 decode_in43
+ decode_in44 decode_in45 decode_in46 decode_in55 decode_in56 decode_in57 decode_in58 decode_in59 decode_in60 decode_in61 decode_in62 OUT3 VDD
+ VDD VSS VSS decode_in8 decode_in9 decode_in10 decode_in11 decode_in12 decode_in13 decode_in14 decode_in15 decode_in24 decode_in25
+ decode_in26 decode_in27 decode_in28 decode_in29 decode_in30 decode_in31 decode_in40 decode_in41 decode_in42 decode_in43 decode_in44
+ decode_in45 decode_in46 decode_in47 decode_in56 decode_in57 decode_in58 decode_in59 decode_in60 decode_in61 decode_in62 or_32
xOut4 decode_in15 decode_in16 decode_in17 decode_in18 decode_in19 decode_in20 decode_in21 decode_in22 decode_in23 decode_in24
+ decode_in25 decode_in26 decode_in27 decode_in28 decode_in29 decode_in30 decode_in47 decode_in48 decode_in49 decode_in50 decode_in51
+ decode_in52 decode_in53 decode_in54 decode_in55 decode_in56 decode_in57 decode_in58 decode_in59 decode_in60 decode_in61 decode_in62 OUT4 VDD
+ VDD VSS VSS decode_in16 decode_in17 decode_in18 decode_in19 decode_in20 decode_in21 decode_in22 decode_in23 decode_in24 decode_in25
+ decode_in26 decode_in27 decode_in28 decode_in29 decode_in30 decode_in31 decode_in48 decode_in49 decode_in50 decode_in51 decode_in52
+ decode_in53 decode_in54 decode_in55 decode_in56 decode_in57 decode_in58 decode_in59 decode_in60 decode_in61 decode_in62 or_32
xOut5 decode_in31 decode_in32 decode_in33 decode_in34 decode_in35 decode_in36 decode_in37 decode_in38 decode_in39 decode_in40
+ decode_in41 decode_in42 decode_in43 decode_in44 decode_in45 decode_in46 decode_in47 decode_in48 decode_in49 decode_in50 decode_in51
+ decode_in52 decode_in53 decode_in54 decode_in55 decode_in56 decode_in57 decode_in58 decode_in59 decode_in60 decode_in61 decode_in62 OUT5 VDD
+ VDD VSS VSS decode_in32 decode_in33 decode_in34 decode_in35 decode_in36 decode_in37 decode_in38 decode_in39 decode_in40 decode_in41
+ decode_in42 decode_in43 decode_in44 decode_in45 decode_in46 decode_in47 decode_in48 decode_in49 decode_in50 decode_in51 decode_in52
+ decode_in53 decode_in54 decode_in55 decode_in56 decode_in57 decode_in58 decode_in59 decode_in60 decode_in61 decode_in62 or_32
.ends


* expanding   symbol:  schematics/comp_top.sym # of pins=6
** sym_path: /home/nwells/xschem/6_bit_flash/schematics/comp_top.sym
** sch_path: /home/nwells/xschem/6_bit_flash/schematics/comp_top.sch
.subckt comp_top VDD vout62 vout61 vout60 vout59 vout58 vout57 vout56 vout55 vout54 vout53 vout52 vout51 vout50 vout49 vout48
+ vout47 vout46 vout45 vout44 vout43 vout42 vout41 vout40 vout39 vout38 vout37 vout36 vout35 vout34 vout33 vout32 vout31 vout30 vout29
+ vout28 vout27 vout26 vout25 vout24 vout23 vout22 vout21 vout20 vout19 vout18 vout17 vout16 vout15 vout14 vout13 vout12 vout11 vout10
+ vout9 vout8 vout7 vout6 vout5 vout4 vout3 vout2 vout1 vout0 VSS vref62 vref61 vref60 vref59 vref58 vref57 vref56 vref55 vref54 vref53
+ vref52 vref51 vref50 vref49 vref48 vref47 vref46 vref45 vref44 vref43 vref42 vref41 vref40 vref39 vref38 vref37 vref36 vref35 vref34
+ vref33 vref32 vref31 vref30 vref29 vref28 vref27 vref26 vref25 vref24 vref23 vref22 vref21 vref20 vref19 vref18 vref17 vref16 vref15
+ vref14 vref13 vref12 vref11 vref10 vref9 vref8 vref7 vref6 vref5 vref4 vref3 vref2 vref1 vref0 VIN clk
*.opin
*+ vout62,vout61,vout60,vout59,vout58,vout57,vout56,vout55,vout54,vout53,vout52,vout51,vout50,vout49,vout48,vout47,vout46,vout45,vout44,vout43,vout42,vout41,vout40,vout39,vout38,vout37,vout36,vout35,vout34,vout33,vout32,vout31,vout30,vout29,vout28,vout27,vout26,vout25,vout24,vout23,vout22,vout21,vout20,vout19,vout18,vout17,vout16,vout15,vout14,vout13,vout12,vout11,vout10,vout9,vout8,vout7,vout6,vout5,vout4,vout3,vout2,vout1,vout0
*.ipin VDD
*.ipin VSS
*.ipin
*+ vref62,vref61,vref60,vref59,vref58,vref57,vref56,vref55,vref54,vref53,vref52,vref51,vref50,vref49,vref48,vref47,vref46,vref45,vref44,vref43,vref42,vref41,vref40,vref39,vref38,vref37,vref36,vref35,vref34,vref33,vref32,vref31,vref30,vref29,vref28,vref27,vref26,vref25,vref24,vref23,vref22,vref21,vref20,vref19,vref18,vref17,vref16,vref15,vref14,vref13,vref12,vref11,vref10,vref9,vref8,vref7,vref6,vref5,vref4,vref3,vref2,vref1,vref0
*.ipin VIN
*.ipin clk
xCOMP62 vout62 VDD VSS VIN vref62 clk comp
xCOMP61 vout61 VDD VSS VIN vref61 clk comp
xCOMP60 vout60 VDD VSS VIN vref60 clk comp
xCOMP59 vout59 VDD VSS VIN vref59 clk comp
xCOMP58 vout58 VDD VSS VIN vref58 clk comp
xCOMP57 vout57 VDD VSS VIN vref57 clk comp
xCOMP56 vout56 VDD VSS VIN vref56 clk comp
xCOMP55 vout55 VDD VSS VIN vref55 clk comp
xCOMP54 vout54 VDD VSS VIN vref54 clk comp
xCOMP53 vout53 VDD VSS VIN vref53 clk comp
xCOMP52 vout52 VDD VSS VIN vref52 clk comp
xCOMP51 vout51 VDD VSS VIN vref51 clk comp
xCOMP50 vout50 VDD VSS VIN vref50 clk comp
xCOMP49 vout49 VDD VSS VIN vref49 clk comp
xCOMP48 vout48 VDD VSS VIN vref48 clk comp
xCOMP47 vout47 VDD VSS VIN vref47 clk comp
xCOMP46 vout46 VDD VSS VIN vref46 clk comp
xCOMP45 vout45 VDD VSS VIN vref45 clk comp
xCOMP44 vout44 VDD VSS VIN vref44 clk comp
xCOMP43 vout43 VDD VSS VIN vref43 clk comp
xCOMP42 vout42 VDD VSS VIN vref42 clk comp
xCOMP41 vout41 VDD VSS VIN vref41 clk comp
xCOMP40 vout40 VDD VSS VIN vref40 clk comp
xCOMP39 vout39 VDD VSS VIN vref39 clk comp
xCOMP38 vout38 VDD VSS VIN vref38 clk comp
xCOMP37 vout37 VDD VSS VIN vref37 clk comp
xCOMP36 vout36 VDD VSS VIN vref36 clk comp
xCOMP35 vout35 VDD VSS VIN vref35 clk comp
xCOMP34 vout34 VDD VSS VIN vref34 clk comp
xCOMP33 vout33 VDD VSS VIN vref33 clk comp
xCOMP32 vout32 VDD VSS VIN vref32 clk comp
xCOMP31 vout31 VDD VSS VIN vref31 clk comp
xCOMP30 vout30 VDD VSS VIN vref30 clk comp
xCOMP29 vout29 VDD VSS VIN vref29 clk comp
xCOMP28 vout28 VDD VSS VIN vref28 clk comp
xCOMP27 vout27 VDD VSS VIN vref27 clk comp
xCOMP26 vout26 VDD VSS VIN vref26 clk comp
xCOMP25 vout25 VDD VSS VIN vref25 clk comp
xCOMP24 vout24 VDD VSS VIN vref24 clk comp
xCOMP23 vout23 VDD VSS VIN vref23 clk comp
xCOMP22 vout22 VDD VSS VIN vref22 clk comp
xCOMP21 vout21 VDD VSS VIN vref21 clk comp
xCOMP20 vout20 VDD VSS VIN vref20 clk comp
xCOMP19 vout19 VDD VSS VIN vref19 clk comp
xCOMP18 vout18 VDD VSS VIN vref18 clk comp
xCOMP17 vout17 VDD VSS VIN vref17 clk comp
xCOMP16 vout16 VDD VSS VIN vref16 clk comp
xCOMP15 vout15 VDD VSS VIN vref15 clk comp
xCOMP14 vout14 VDD VSS VIN vref14 clk comp
xCOMP13 vout13 VDD VSS VIN vref13 clk comp
xCOMP12 vout12 VDD VSS VIN vref12 clk comp
xCOMP11 vout11 VDD VSS VIN vref11 clk comp
xCOMP10 vout10 VDD VSS VIN vref10 clk comp
xCOMP9 vout9 VDD VSS VIN vref9 clk comp
xCOMP8 vout8 VDD VSS VIN vref8 clk comp
xCOMP7 vout7 VDD VSS VIN vref7 clk comp
xCOMP6 vout6 VDD VSS VIN vref6 clk comp
xCOMP5 vout5 VDD VSS VIN vref5 clk comp
xCOMP4 vout4 VDD VSS VIN vref4 clk comp
xCOMP3 vout3 VDD VSS VIN vref3 clk comp
xCOMP2 vout2 VDD VSS VIN vref2 clk comp
xCOMP1 vout1 VDD VSS VIN vref1 clk comp
xCOMP0 vout0 VDD VSS VIN vref0 clk comp
.ends


* expanding   symbol:  schematics/ideal_comp.sym # of pins=5
** sym_path: /home/nwells/xschem/6_bit_flash/schematics/ideal_comp.sym
** sch_path: /home/nwells/xschem/6_bit_flash/schematics/ideal_comp.sch
.subckt ideal_comp vdd vss vinp vout vinn  bw=100Meg gain=100 vcmh=1.6 vcml=0.2 vios=50m
*.ipin vdd
*.opin vout
*.ipin vss
*.ipin vinp
*.ipin vinn
B1 vp vss V = {V(vinp)<vcmh ? (V(vinp) < vcml ? vcml: V(vinp)) : vcmh} m=1
B2 vn vss V = {V(vinn)<vcmh ? (V(vinn) < vcml ? vcml: V(vinn) + vios) : vcmh} m=1
B3 net1 vss V = {gain*(V(vp)-V(vn)) < V(vdd) ? (gain*(V(vp)-V(vn)) < V(vss) ? V(vss) : (gain*(V(vp)-V(vn)))) : V(vdd)} m=1
R1 vout net1 {1/(2*3.1415*bw*1p)} m=1
C1 vout vss 1p m=1
.ends


* expanding   symbol:  schematics/or_32.sym # of pins=68
** sym_path: /home/nwells/xschem/6_bit_flash/schematics/or_32.sym
** sch_path: /home/nwells/xschem/6_bit_flash/schematics/or_32.sch
.subckt or_32 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 I16 I17 I18 I19 I20 I21 I22 I23 I24 I25 I26 I27 I28 I29 I30 I31
+ I32 O VPWR VPB VGND VNB I1_AND I2_AND I3_AND I4_AND I5_AND I6_AND I7_AND I8_AND I9_AND I10_AND I11_AND I12_AND I13_AND I14_AND
+ I15_AND I16_AND I17_AND I18_AND I19_AND I20_AND I21_AND I22_AND I23_AND I24_AND I25_AND I26_AND I27_AND I28_AND I29_AND I30_AND I31_AND
*.ipin I1
*.ipin I2
*.ipin I12
*.ipin I3
*.ipin I4
*.ipin I5
*.ipin I6
*.ipin I7
*.ipin I8
*.ipin I9
*.ipin I10
*.ipin I11
*.ipin I13
*.ipin I14
*.ipin I15
*.ipin I16
*.ipin I17
*.ipin I18
*.ipin I19
*.ipin I20
*.ipin I21
*.ipin I22
*.ipin I23
*.ipin I24
*.ipin I25
*.ipin I26
*.ipin I27
*.ipin I28
*.ipin I29
*.ipin I30
*.ipin I31
*.ipin I32
*.opin O
*.ipin VGND
*.ipin VNB
*.ipin VPB
*.ipin VPWR
*.ipin I1_AND
*.ipin I2_AND
*.ipin I12_AND
*.ipin I3_AND
*.ipin I4_AND
*.ipin I5_AND
*.ipin I6_AND
*.ipin I7_AND
*.ipin I8_AND
*.ipin I9_AND
*.ipin I10_AND
*.ipin I11_AND
*.ipin I13_AND
*.ipin I14_AND
*.ipin I15_AND
*.ipin I16_AND
*.ipin I17_AND
*.ipin I18_AND
*.ipin I19_AND
*.ipin I20_AND
*.ipin I21_AND
*.ipin I22_AND
*.ipin I23_AND
*.ipin I24_AND
*.ipin I25_AND
*.ipin I26_AND
*.ipin I27_AND
*.ipin I28_AND
*.ipin I29_AND
*.ipin I30_AND
*.ipin I31_AND
x10 net3 net4 net5 net6 VGND VNB VPB VPWR net1 sky130_fd_sc_hd__or4_1
x9 net1 net2 VGND VNB VPB VPWR O sky130_fd_sc_hd__or2_0
x1 I1 I1_AND I2 I2_AND I3 I3_AND I4 I4_AND VPWR VPB VGND VNB net3 or_4_and_2
x2 I5 I5_AND I6 I6_AND I7 I7_AND I8 I8_AND VPWR VPB VGND VNB net4 or_4_and_2
x3 I9 I9_AND I10 I10_AND I11 I11_AND I12 I12_AND VPWR VPB VGND VNB net5 or_4_and_2
x4 I13 I13_AND I14 I14_AND I15 I15_AND I16 I16_AND VPWR VPB VGND VNB net6 or_4_and_2
x5 net7 net8 net9 net10 VGND VNB VPB VPWR net2 sky130_fd_sc_hd__or4_1
x6 I17 I17_AND I18 I18_AND I19 I19_AND I20 I20_AND VPWR VPB VGND VNB net7 or_4_and_2
x7 I21 I21_AND I22 I22_AND I23 I23_AND I24 I24_AND VPWR VPB VGND VNB net8 or_4_and_2
x8 I25 I25_AND I26 I26_AND I27 I27_AND I28 I28_AND VPWR VPB VGND VNB net9 or_4_and_2
x11 I29 I29_AND I30 I30_AND I31 I31_AND I32 VGND VPWR VPB VGND VNB net10 or_4_and_2
.ends


* expanding   symbol:  schematics/comp.sym # of pins=6
** sym_path: /home/nwells/xschem/6_bit_flash/schematics/comp.sym
** sch_path: /home/nwells/xschem/6_bit_flash/schematics/comp.sch
.subckt comp vout vdd vss vinp vinn clk
*.ipin vdd
*.opin vout
*.ipin vss
*.ipin vinp
*.ipin vinn
*.ipin clk
XM1 vinp_d vinp vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM2 vinn_d vinn vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM3 voutn voutp vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=7.5 nf=1 ad=2.175 as=2.175 pd=15.58 ps=15.58 nrd=0.0386666666666667
+ nrs=0.0386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM4 voutp voutn vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=7.5 nf=1 ad=2.175 as=2.175 pd=15.58 ps=15.58 nrd=0.0386666666666667
+ nrs=0.0386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM5 vinp_d vinn_d vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=7.5 nf=1 ad=2.175 as=2.175 pd=15.58 ps=15.58 nrd=0.0386666666666667
+ nrs=0.0386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM6 vinn_d vinp_d vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=7.5 nf=1 ad=2.175 as=2.175 pd=15.58 ps=15.58 nrd=0.0386666666666667
+ nrs=0.0386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM7 voutn clk vinp_d vss sky130_fd_pr__nfet_01v8 L=0.18 W=1.5 nf=1 ad=0.435 as=0.435 pd=3.58 ps=3.58 nrd=0.193333333333333
+ nrs=0.193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM8 voutp clk vinn_d vss sky130_fd_pr__nfet_01v8 L=0.18 W=1.5 nf=1 ad=0.435 as=0.435 pd=3.58 ps=3.58 nrd=0.193333333333333
+ nrs=0.193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM9 voutn clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=4 nf=1 ad=1.16 as=1.16 pd=8.58 ps=8.58 nrd=0.0725 nrs=0.0725 sa=0 sb=0 sd=0
+ mult=1 m=1
XM10 voutp clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=4 nf=1 ad=1.16 as=1.16 pd=8.58 ps=8.58 nrd=0.0725 nrs=0.0725 sa=0 sb=0
+ sd=0 mult=1 m=1
xBUFF voutp vss vss vdd vdd voutp_buff sky130_fd_sc_hd__buf_6
xBUFF1 voutn vss vss vdd vdd voutn_buff sky130_fd_sc_hd__buf_6
I0 pa_m1_s vss 10u
XM11 v_m1_d voutp_buff pa_m1_s vss sky130_fd_pr__nfet_01v8 L=0.15 W=50 nf=1 ad=14.5 as=14.5 pd=100.58 ps=100.58 nrd=0.0058
+ nrs=0.0058 sa=0 sb=0 sd=0 mult=1 m=1
XM12 vout voutn_buff pa_m1_s vss sky130_fd_pr__nfet_01v8 L=0.15 W=50 nf=1 ad=14.5 as=14.5 pd=100.58 ps=100.58 nrd=0.0058
+ nrs=0.0058 sa=0 sb=0 sd=0 mult=1 m=1
XM13 v_m1_d v_m1_d vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0
+ sd=0 mult=1 m=1
XM14 vout v_m1_d vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
.ends


* expanding   symbol:  schematics/or_4_and_2.sym # of pins=13
** sym_path: /home/nwells/xschem/6_bit_flash/schematics/or_4_and_2.sym
** sch_path: /home/nwells/xschem/6_bit_flash/schematics/or_4_and_2.sch
.subckt or_4_and_2 I1 I1_AND I2 I2_AND I3 I3_AND I4 I4_AND VPWR VPB VGND VNB O
*.opin O
*.ipin I1
*.ipin I2
*.ipin I3
*.ipin I4
*.ipin I1_AND
*.ipin I2_AND
*.ipin I3_AND
*.ipin I4_AND
*.ipin VGND
*.ipin VNB
*.ipin VPB
*.ipin VPWR
x1 net3 net1 net4 net2 VGND VNB VPB VPWR O sky130_fd_sc_hd__or4_1
x2 I2 net5 VGND VNB VPB VPWR net1 sky130_fd_sc_hd__and2_0
x3 I1 net6 VGND VNB VPB VPWR net3 sky130_fd_sc_hd__and2_0
x4 I4 net7 VGND VNB VPB VPWR net2 sky130_fd_sc_hd__and2_0
x5 I3 net8 VGND VNB VPB VPWR net4 sky130_fd_sc_hd__and2_0
x6 I2_AND VGND VNB VPB VPWR net5 sky130_fd_sc_hd__inv_1
x7 I1_AND VGND VNB VPB VPWR net6 sky130_fd_sc_hd__inv_1
x8 I3_AND VGND VNB VPB VPWR net8 sky130_fd_sc_hd__inv_1
x9 I4_AND VGND VNB VPB VPWR net7 sky130_fd_sc_hd__inv_1
.ends

**** begin user architecture code

.subckt decoder_6bit_cell vdd out5 out4 out3 out2 out1 out0 dec_in62 dec_in61 dec_in60 dec_in59 dec_in58 dec_in57 dec_in56 dec_in55 dec_in54 dec_in53 dec_in52 dec_in51 dec_in50 dec_in49 dec_in48 dec_in47 dec_in46 dec_in45 dec_in44 dec_in43 dec_in42 dec_in41 dec_in40 dec_in39 dec_in38 dec_in37 dec_in36 dec_in35 dec_in34 dec_in33 dec_in32 dec_in31 dec_in30 dec_in29 dec_in28 dec_in27 dec_in26 dec_in25 dec_in24 dec_in23 dec_in22 dec_in21 dec_in20 dec_in19 dec_in18 dec_in17 dec_in16 dec_in15 dec_in14 dec_in13 dec_in12 dec_in11 dec_in10 dec_in9 dec_in8 dec_in7 dec_in6 dec_in5 dec_in4 dec_in3 dec_in2 dec_in1 dec_in0 vss vref
N1 vdd out5 out4 out3 out2 out1 out0 dec_in62 dec_in61 dec_in60 dec_in59 dec_in58 dec_in57 dec_in56 dec_in55 dec_in54 dec_in53 dec_in52 dec_in51 dec_in50 dec_in49 dec_in48 dec_in47 dec_in46 dec_in45 dec_in44 dec_in43 dec_in42 dec_in41 dec_in40 dec_in39 dec_in38 dec_in37 dec_in36 dec_in35 dec_in34 dec_in33 dec_in32 dec_in31 dec_in30 dec_in29 dec_in28 dec_in27 dec_in26 dec_in25 dec_in24 dec_in23 dec_in22 dec_in21 dec_in20 dec_in19 dec_in18 dec_in17 dec_in16 dec_in15 dec_in14 dec_in13 dec_in12 dec_in11 dec_in10 dec_in9 dec_in8 dec_in7 dec_in6 dec_in5 dec_in4 dec_in3 dec_in2 dec_in1 dec_in0 vss vref decoder_6bit_model
.ends decoder_6bit_cell

.model decoder_6bit_model decoder_6bit



.control
* following line specifies the location for the .osdi file so ngspice can use it.
* working dir set in tcl in startup script as pwd in top location
pre_osdi /home/nwells/xschem/6_bit_flash/schematics/verilog_a/ideal_decoder.osdi
.endc


.subckt ideal_comp_cell VDD VSS INP INN VOUT
N1 vdd vss inp inn vout ideal_comp_model
.ends ideal_comp_cell

.model ideal_comp_model ideal_comp


.control
* following line specifies the location for the .osdi file so ngspice can use it.
* working dir set in tcl in startup script as pwd in top location
pre_osdi /home/nwells/xschem/6_bit_flash/schematics/verilog_a/ideal_comp.osdi
.endc

**** end user architecture code
.end
