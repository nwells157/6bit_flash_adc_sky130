** sch_path: /home/nwells/xschem/6_bit_flash/schematics/adc_top.sch
**.subckt adc_top OUT5,OUT4,OUT3,OUT2,OUT1,OUT0 VDD
*+ vref62,vref61,vref60,vref59,vref58,vref57,vref56,vref55,vref54,vref53,vref52,vref51,vref50,vref49,vref48,vref47,vref46,vref45,vref44,vref43,vref42,vref41,vref40,vref39,vref38,vref37,vref36,vref35,vref34,vref33,vref32,vref31,vref30,vref29,vref28,vref27,vref26,vref25,vref24,vref23,vref22,vref21,vref20,vref19,vref18,vref17,vref16,vref15,vref14,vref13,vref12,vref11,vref10,vref9,vref8,vref7,vref6,vref5,vref4,vref3,vref2,vref1,vref0 VSS
*+ comp_out62,comp_out61,comp_out60,comp_out59,comp_out58,comp_out57,comp_out56,comp_out55,comp_out54,comp_out53,comp_out52,comp_out51,comp_out50,comp_out49,comp_out48,comp_out47,comp_out46,comp_out45,comp_out44,comp_out43,comp_out42,comp_out41,comp_out40,comp_out39,comp_out38,comp_out37,comp_out36,comp_out35,comp_out34,comp_out33,comp_out32,comp_out31,comp_out30,comp_out29,comp_out28,comp_out27,comp_out26,comp_out25,comp_out24,comp_out23,comp_out22,comp_out21,comp_out20,comp_out19,comp_out18,comp_out17,comp_out16,comp_out15,comp_out14,comp_out13,comp_out12,comp_out11,comp_out10,comp_out9,comp_out8,comp_out7,comp_out6,comp_out5,comp_out4,comp_out3,comp_out2,comp_out1,comp_out0 VIN VREF clk
*.ipin VDD
*.ipin VSS
*.ipin VIN
*.ipin VREF
*.opin OUT5,OUT4,OUT3,OUT2,OUT1,OUT0
*.iopin
*+ vref62,vref61,vref60,vref59,vref58,vref57,vref56,vref55,vref54,vref53,vref52,vref51,vref50,vref49,vref48,vref47,vref46,vref45,vref44,vref43,vref42,vref41,vref40,vref39,vref38,vref37,vref36,vref35,vref34,vref33,vref32,vref31,vref30,vref29,vref28,vref27,vref26,vref25,vref24,vref23,vref22,vref21,vref20,vref19,vref18,vref17,vref16,vref15,vref14,vref13,vref12,vref11,vref10,vref9,vref8,vref7,vref6,vref5,vref4,vref3,vref2,vref1,vref0
*.iopin
*+ comp_out62,comp_out61,comp_out60,comp_out59,comp_out58,comp_out57,comp_out56,comp_out55,comp_out54,comp_out53,comp_out52,comp_out51,comp_out50,comp_out49,comp_out48,comp_out47,comp_out46,comp_out45,comp_out44,comp_out43,comp_out42,comp_out41,comp_out40,comp_out39,comp_out38,comp_out37,comp_out36,comp_out35,comp_out34,comp_out33,comp_out32,comp_out31,comp_out30,comp_out29,comp_out28,comp_out27,comp_out26,comp_out25,comp_out24,comp_out23,comp_out22,comp_out21,comp_out20,comp_out19,comp_out18,comp_out17,comp_out16,comp_out15,comp_out14,comp_out13,comp_out12,comp_out11,comp_out10,comp_out9,comp_out8,comp_out7,comp_out6,comp_out5,comp_out4,comp_out3,comp_out2,comp_out1,comp_out0
*.ipin clk
xREF_LADDER VDD vref62 vref61 vref60 vref59 vref58 vref57 vref56 vref55 vref54 vref53 vref52 vref51 vref50 vref49 vref48 vref47
+ vref46 vref45 vref44 vref43 vref42 vref41 vref40 vref39 vref38 vref37 vref36 vref35 vref34 vref33 vref32 vref31 vref30 vref29 vref28
+ vref27 vref26 vref25 vref24 vref23 vref22 vref21 vref20 vref19 vref18 vref17 vref16 vref15 vref14 vref13 vref12 vref11 vref10 vref9
+ vref8 vref7 vref6 vref5 vref4 vref3 vref2 vref1 vref0 VSS ref_ladder_top
xVERILOGA_DECODER_TOP VDD OUT5 OUT4 OUT3 OUT2 OUT1 OUT0 comp_out62 comp_out61 comp_out60 comp_out59 comp_out58 comp_out57
+ comp_out56 comp_out55 comp_out54 comp_out53 comp_out52 comp_out51 comp_out50 comp_out49 comp_out48 comp_out47 comp_out46 comp_out45
+ comp_out44 comp_out43 comp_out42 comp_out41 comp_out40 comp_out39 comp_out38 comp_out37 comp_out36 comp_out35 comp_out34 comp_out33
+ comp_out32 comp_out31 comp_out30 comp_out29 comp_out28 comp_out27 comp_out26 comp_out25 comp_out24 comp_out23 comp_out22 comp_out21
+ comp_out20 comp_out19 comp_out18 comp_out17 comp_out16 comp_out15 comp_out14 comp_out13 comp_out12 comp_out11 comp_out10 comp_out9 comp_out8
+ comp_out7 comp_out6 comp_out5 comp_out4 comp_out3 comp_out2 comp_out1 comp_out0 VSS VREF decoder_6bit_cell
xIDEAL_COMP_TOP comp_out62 comp_out61 comp_out60 comp_out59 comp_out58 comp_out57 comp_out56 comp_out55 comp_out54 comp_out53
+ comp_out52 comp_out51 comp_out50 comp_out49 comp_out48 comp_out47 comp_out46 comp_out45 comp_out44 comp_out43 comp_out42 comp_out41
+ comp_out40 comp_out39 comp_out38 comp_out37 comp_out36 comp_out35 comp_out34 comp_out33 comp_out32 comp_out31 comp_out30 comp_out29
+ comp_out28 comp_out27 comp_out26 comp_out25 comp_out24 comp_out23 comp_out22 comp_out21 comp_out20 comp_out19 comp_out18 comp_out17
+ comp_out16 comp_out15 comp_out14 comp_out13 comp_out12 comp_out11 comp_out10 comp_out9 comp_out8 comp_out7 comp_out6 comp_out5 comp_out4
+ comp_out3 comp_out2 comp_out1 comp_out0 VDD VSS vref62 vref61 vref60 vref59 vref58 vref57 vref56 vref55 vref54 vref53 vref52 vref51 vref50
+ vref49 vref48 vref47 vref46 vref45 vref44 vref43 vref42 vref41 vref40 vref39 vref38 vref37 vref36 vref35 vref34 vref33 vref32 vref31
+ vref30 vref29 vref28 vref27 vref26 vref25 vref24 vref23 vref22 vref21 vref20 vref19 vref18 vref17 vref16 vref15 vref14 vref13 vref12
+ vref11 vref10 vref9 vref8 vref7 vref6 vref5 vref4 vref3 vref2 vref1 vref0 VIN comp_top_ideal
**.ends
**** begin user architecture code

.subckt decoder_6bit_cell vdd out5 out4 out3 out2 out1 out0 dec_in62 dec_in61 dec_in60 dec_in59 dec_in58 dec_in57 dec_in56 dec_in55 dec_in54 dec_in53 dec_in52 dec_in51 dec_in50 dec_in49 dec_in48 dec_in47 dec_in46 dec_in45 dec_in44 dec_in43 dec_in42 dec_in41 dec_in40 dec_in39 dec_in38 dec_in37 dec_in36 dec_in35 dec_in34 dec_in33 dec_in32 dec_in31 dec_in30 dec_in29 dec_in28 dec_in27 dec_in26 dec_in25 dec_in24 dec_in23 dec_in22 dec_in21 dec_in20 dec_in19 dec_in18 dec_in17 dec_in16 dec_in15 dec_in14 dec_in13 dec_in12 dec_in11 dec_in10 dec_in9 dec_in8 dec_in7 dec_in6 dec_in5 dec_in4 dec_in3 dec_in2 dec_in1 dec_in0 vss vref
N1 vdd out5 out4 out3 out2 out1 out0 dec_in62 dec_in61 dec_in60 dec_in59 dec_in58 dec_in57 dec_in56 dec_in55 dec_in54 dec_in53 dec_in52 dec_in51 dec_in50 dec_in49 dec_in48 dec_in47 dec_in46 dec_in45 dec_in44 dec_in43 dec_in42 dec_in41 dec_in40 dec_in39 dec_in38 dec_in37 dec_in36 dec_in35 dec_in34 dec_in33 dec_in32 dec_in31 dec_in30 dec_in29 dec_in28 dec_in27 dec_in26 dec_in25 dec_in24 dec_in23 dec_in22 dec_in21 dec_in20 dec_in19 dec_in18 dec_in17 dec_in16 dec_in15 dec_in14 dec_in13 dec_in12 dec_in11 dec_in10 dec_in9 dec_in8 dec_in7 dec_in6 dec_in5 dec_in4 dec_in3 dec_in2 dec_in1 dec_in0 vss vref decoder_6bit_model
.ends decoder_6bit_cell

.model decoder_6bit_model decoder_6bit



.control
* following line specifies the location for the .osdi file so ngspice can use it.
* working dir set in tcl in startup script as pwd in top location
pre_osdi /home/nwells/xschem/6_bit_flash/schematics/verilog_a/ideal_decoder.osdi
.endc

**** end user architecture code
.end
