** sch_path: /home/nwells/xschem/6_bit_flash/schematics/comp.sch
**.subckt comp pa_voutp vdd vout pa_voutn vss vinp latch_voutp latch_voutn vinn pa_m1_s
*.ipin vdd
*.opin vout
*.ipin vss
*.ipin vinp
*.ipin vinn
*.iopin pa_voutp
*.iopin pa_voutn
*.iopin latch_voutp
*.iopin latch_voutn
*.iopin pa_m1_s
I0 pa_m1_s vss 10u
XM1 v_m1_d vinp pa_m1_s pa_m1_s sky130_fd_pr__nfet_01v8 L=0.5 W=20 nf=1 ad=5.8 as=5.8 pd=40.58 ps=40.58 nrd=0.0145 nrs=0.0145 sa=0
+ sb=0 sd=0 mult=1 m=1
XM2 net1 vinn pa_m1_s pa_m1_s sky130_fd_pr__nfet_01v8 L=0.5 W=20 nf=1 ad=5.8 as=5.8 pd=40.58 ps=40.58 nrd=0.0145 nrs=0.0145 sa=0
+ sb=0 sd=0 mult=1 m=1
XM3 v_m1_d v_m1_d vdd vdd sky130_fd_pr__pfet_01v8 L=2 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
XM4 net1 v_m1_d vdd vdd sky130_fd_pr__pfet_01v8 L=2 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
XM5 net2 net1 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM6 net2 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
XM7 vout net2 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM8 vout net2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
**.ends
.end
