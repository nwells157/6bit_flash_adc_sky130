** IDEAL_DAC_TEMP flat netlist
.end
